module FSM(
  input In1,
  input RST,
  input CLK, 
  output reg Out1
);
