// ProjectSystem.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module ProjectSystem (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule
