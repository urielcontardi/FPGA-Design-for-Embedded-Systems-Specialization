// Embed.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Embed (
		input  wire        altpll_1_areset_conduit_export,      //      altpll_1_areset_conduit.export
		output wire        altpll_1_locked_conduit_export,      //      altpll_1_locked_conduit.export
		input  wire        clk_clk,                             //                          clk.clk
		input  wire        clk_0_clk,                           //                        clk_0.clk
		output wire [12:0] dram_addr,                           //                         dram.addr
		output wire [1:0]  dram_ba,                             //                             .ba
		output wire        dram_cas_n,                          //                             .cas_n
		output wire        dram_cke,                            //                             .cke
		output wire        dram_cs_n,                           //                             .cs_n
		inout  wire [15:0] dram_dq,                             //                             .dq
		output wire [1:0]  dram_dqm,                            //                             .dqm
		output wire        dram_ras_n,                          //                             .ras_n
		output wire        dram_we_n,                           //                             .we_n
		output wire        dram_clk_clk,                        //                     dram_clk.clk
		input  wire        gsensor_MISO,                        //                      gsensor.MISO
		output wire        gsensor_MOSI,                        //                             .MOSI
		output wire        gsensor_SCLK,                        //                             .SCLK
		output wire        gsensor_SS_n,                        //                             .SS_n
		output wire [9:0]  ledr_export,                         //                         ledr.export
		input  wire        modular_adc_0_adc_pll_locked_export, // modular_adc_0_adc_pll_locked.export
		input  wire        reset_reset_n,                       //                        reset.reset_n
		input  wire        reset_0_reset_n,                     //                      reset_0.reset_n
		input  wire [9:0]  sw_export                            //                           sw.export
	);

	wire         altpll_1_c0_clk;                                               // altpll_1:c0 -> modular_adc_0:adc_pll_clock_clk
	wire         altpll_0_c0_clk;                                               // altpll_0:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, mm_clock_crossing_bridge_0:s0_clk, mm_interconnect_0:altpll_0_c0_clk, nios2_gen2_0:clk, onchip_flash_0:clock, onchip_memory2_0:clk, rst_controller_004:clk, sdram:clk, spi_0:clk]
	wire         altpll_0_c2_clk;                                               // altpll_0:c2 -> [irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, jtag_uart_0:clk, led_pio:clk, mm_clock_crossing_bridge_0:m0_clk, mm_interconnect_1:altpll_0_c2_clk, rst_controller_002:clk, slide_pio:clk, sysid:clock, timer_0:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                             // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                          // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                          // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                              // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                           // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                 // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                        // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                            // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] master_0_master_readdata;                                      // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                                   // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                       // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                          // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                    // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                                 // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                         // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                     // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                      // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                   // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                       // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                          // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_readdata;                 // onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	wire   [0:0] mm_interconnect_0_onchip_flash_0_csr_address;                  // mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	wire         mm_interconnect_0_onchip_flash_0_csr_read;                     // mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	wire         mm_interconnect_0_onchip_flash_0_csr_write;                    // mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_csr_writedata;                // mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_readdata;                // onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	wire         mm_interconnect_0_onchip_flash_0_data_waitrequest;             // onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	wire  [18:0] mm_interconnect_0_onchip_flash_0_data_address;                 // mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	wire         mm_interconnect_0_onchip_flash_0_data_read;                    // mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	wire         mm_interconnect_0_onchip_flash_0_data_readdatavalid;           // onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	wire         mm_interconnect_0_onchip_flash_0_data_write;                   // mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	wire  [31:0] mm_interconnect_0_onchip_flash_0_data_writedata;               // mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	wire   [3:0] mm_interconnect_0_onchip_flash_0_data_burstcount;              // mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;       // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;    // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata;      // mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest;   // mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid; // mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;              // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                 // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;              // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                   // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;               // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                   // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                         // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                           // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                        // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                            // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                               // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                         // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                      // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                              // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                          // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_modular_adc_0_sample_store_csr_readdata;     // modular_adc_0:sample_store_csr_readdata -> mm_interconnect_0:modular_adc_0_sample_store_csr_readdata
	wire   [6:0] mm_interconnect_0_modular_adc_0_sample_store_csr_address;      // mm_interconnect_0:modular_adc_0_sample_store_csr_address -> modular_adc_0:sample_store_csr_address
	wire         mm_interconnect_0_modular_adc_0_sample_store_csr_read;         // mm_interconnect_0:modular_adc_0_sample_store_csr_read -> modular_adc_0:sample_store_csr_read
	wire         mm_interconnect_0_modular_adc_0_sample_store_csr_write;        // mm_interconnect_0:modular_adc_0_sample_store_csr_write -> modular_adc_0:sample_store_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_0_sample_store_csr_writedata;    // mm_interconnect_0:modular_adc_0_sample_store_csr_writedata -> modular_adc_0:sample_store_csr_writedata
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_readdata;        // modular_adc_0:sequencer_csr_readdata -> mm_interconnect_0:modular_adc_0_sequencer_csr_readdata
	wire   [0:0] mm_interconnect_0_modular_adc_0_sequencer_csr_address;         // mm_interconnect_0:modular_adc_0_sequencer_csr_address -> modular_adc_0:sequencer_csr_address
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_read;            // mm_interconnect_0:modular_adc_0_sequencer_csr_read -> modular_adc_0:sequencer_csr_read
	wire         mm_interconnect_0_modular_adc_0_sequencer_csr_write;           // mm_interconnect_0:modular_adc_0_sequencer_csr_write -> modular_adc_0:sequencer_csr_write
	wire  [31:0] mm_interconnect_0_modular_adc_0_sequencer_csr_writedata;       // mm_interconnect_0:modular_adc_0_sequencer_csr_writedata -> modular_adc_0:sequencer_csr_writedata
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;           // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_readdata;             // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;              // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;                 // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;                // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_writedata;            // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                 // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                  // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                     // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                    // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_0_altpll_1_pll_slave_readdata;                 // altpll_1:readdata -> mm_interconnect_0:altpll_1_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_1_pll_slave_address;                  // mm_interconnect_0:altpll_1_pll_slave_address -> altpll_1:address
	wire         mm_interconnect_0_altpll_1_pll_slave_read;                     // mm_interconnect_0:altpll_1_pll_slave_read -> altpll_1:read
	wire         mm_interconnect_0_altpll_1_pll_slave_write;                    // mm_interconnect_0:altpll_1_pll_slave_write -> altpll_1:write
	wire  [31:0] mm_interconnect_0_altpll_1_pll_slave_writedata;                // mm_interconnect_0:altpll_1_pll_slave_writedata -> altpll_1:writedata
	wire         mm_clock_crossing_bridge_0_m0_waitrequest;                     // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_0_m0_readdata;                        // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire         mm_clock_crossing_bridge_0_m0_debugaccess;                     // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_0_m0_address;                         // mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_address
	wire         mm_clock_crossing_bridge_0_m0_read;                            // mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_read
	wire   [3:0] mm_clock_crossing_bridge_0_m0_byteenable;                      // mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_byteenable
	wire         mm_clock_crossing_bridge_0_m0_readdatavalid;                   // mm_interconnect_1:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_0_m0_writedata;                       // mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_writedata
	wire         mm_clock_crossing_bridge_0_m0_write;                           // mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_write
	wire   [0:0] mm_clock_crossing_bridge_0_m0_burstcount;                      // mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_0_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;    // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;      // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest;   // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;       // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;          // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;         // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;     // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                 // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_led_pio_s1_chipselect;                       // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;                         // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                          // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                            // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;                        // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_1_slide_pio_s1_chipselect;                     // mm_interconnect_1:slide_pio_s1_chipselect -> slide_pio:chipselect
	wire  [31:0] mm_interconnect_1_slide_pio_s1_readdata;                       // slide_pio:readdata -> mm_interconnect_1:slide_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_slide_pio_s1_address;                        // mm_interconnect_1:slide_pio_s1_address -> slide_pio:address
	wire         mm_interconnect_1_slide_pio_s1_write;                          // mm_interconnect_1:slide_pio_s1_write -> slide_pio:write_n
	wire  [31:0] mm_interconnect_1_slide_pio_s1_writedata;                      // mm_interconnect_1:slide_pio_s1_writedata -> slide_pio:writedata
	wire         mm_interconnect_1_timer_0_s1_chipselect;                       // mm_interconnect_1:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_1_timer_0_s1_readdata;                         // timer_0:readdata -> mm_interconnect_1:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_0_s1_address;                          // mm_interconnect_1:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_1_timer_0_s1_write;                            // mm_interconnect_1:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_1_timer_0_s1_writedata;                        // mm_interconnect_1:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                                      // spi_0:irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                          // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver1_irq;                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                 // slide_pio:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                      // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                             // timer_0:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver3_irq;                                      // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                             // jtag_uart_0:av_irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver4_irq;                                      // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                             // modular_adc_0:sample_store_irq_irq -> irq_synchronizer_003:receiver_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         nios2_gen2_0_debug_reset_request_reset;                        // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2, rst_controller_004:reset_in2]
	wire         master_0_master_reset_reset;                                   // master_0:master_reset_reset -> [rst_controller:reset_in3, rst_controller_001:reset_in3, rst_controller_002:reset_in3, rst_controller_003:reset_in3, rst_controller_004:reset_in3]
	wire         rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [altpll_1:reset, irq_synchronizer_003:receiver_reset, mm_interconnect_0:master_0_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:modular_adc_0_reset_sink_reset_bridge_in_reset_reset, modular_adc_0:reset_sink_reset_n]
	wire         rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> [irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, jtag_uart_0:rst_n, led_pio:reset_n, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset, slide_pio:reset_n, sysid:reset_n, timer_0:reset_n]
	wire         rst_controller_003_reset_out_reset;                            // rst_controller_003:reset_out -> master_0:clk_reset_reset
	wire         rst_controller_004_reset_out_reset;                            // rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_flash_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram:reset_n, spi_0:reset_n]
	wire         rst_controller_004_reset_out_reset_req;                        // rst_controller_004:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	Embed_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (dram_clk_clk),                                   //                    c1.clk
		.c2                 (altpll_0_c2_clk),                                //                    c2.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	Embed_altpll_1 altpll_1 (
		.clk                (clk_0_clk),                                      //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_1_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_1_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_1_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_1_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_1_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_1_c0_clk),                                //                    c0.clk
		.areset             (altpll_1_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_1_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c1                 (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	Embed_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c2_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_002_receiver_irq)                            //               irq.irq
	);

	Embed_led_pio led_pio (
		.clk        (altpll_0_c2_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),   //                    .readdata
		.out_port   (ledr_export)                              // external_connection.export
	);

	Embed_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_0_clk),                          //          clk.clk
		.clk_reset_reset      (rst_controller_003_reset_out_reset), //    clk_reset.reset
		.master_address       (master_0_master_address),            //       master.address
		.master_readdata      (master_0_master_readdata),           //             .readdata
		.master_read          (master_0_master_read),               //             .read
		.master_write         (master_0_master_write),              //             .write
		.master_writedata     (master_0_master_writedata),          //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),        //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid),      //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),         //             .byteenable
		.master_reset_reset   (master_0_master_reset_reset)         // master_reset.reset
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (altpll_0_c2_clk),                                               //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (altpll_0_c0_clk),                                               //   s0_clk.clk
		.s0_reset         (rst_controller_004_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)                      //         .debugaccess
	);

	Embed_modular_adc_0 #(
		.is_this_first_or_second_adc (1)
	) modular_adc_0 (
		.clock_clk                  (clk_0_clk),                                                  //            clock.clk
		.reset_sink_reset_n         (~rst_controller_001_reset_out_reset),                        //       reset_sink.reset_n
		.adc_pll_clock_clk          (altpll_1_c0_clk),                                            //    adc_pll_clock.clk
		.adc_pll_locked_export      (modular_adc_0_adc_pll_locked_export),                        //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_0_modular_adc_0_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_0_modular_adc_0_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_0_modular_adc_0_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_0_modular_adc_0_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_0_modular_adc_0_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_0_modular_adc_0_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_0_modular_adc_0_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_0_modular_adc_0_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       (irq_synchronizer_003_receiver_irq)                           // sample_store_irq.irq
	);

	Embed_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c0_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_004_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_004_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       (""),
		.INIT_FILENAME_SIM                   (""),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M50DAF484C6GES"),
		.DEVICE_ID                           ("50"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (8191),
		.SECTOR2_START_ADDR                  (8192),
		.SECTOR2_END_ADDR                    (16383),
		.SECTOR3_START_ADDR                  (16384),
		.SECTOR3_END_ADDR                    (114687),
		.SECTOR4_START_ADDR                  (114688),
		.SECTOR4_END_ADDR                    (188415),
		.SECTOR5_START_ADDR                  (188416),
		.SECTOR5_END_ADDR                    (360447),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (360447),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (16383),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (3),
		.SECTOR4_MAP                         (4),
		.SECTOR5_MAP                         (5),
		.ADDR_RANGE1_END_ADDR                (360447),
		.ADDR_RANGE2_END_ADDR                (360447),
		.ADDR_RANGE1_OFFSET                  (2048),
		.ADDR_RANGE2_OFFSET                  (0),
		.ADDR_RANGE3_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (19),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (4),
		.SECTOR_READ_PROTECTION_MODE         (28),
		.FLASH_SEQ_READ_DATA_COUNT           (4),
		.FLASH_ADDR_ALIGNMENT_BITS           (2),
		.FLASH_READ_CYCLE_MAX_INDEX          (5),
		.FLASH_RESET_CYCLE_MAX_INDEX         (20),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (96),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (28000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (24400),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (1),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("False"),
		.IS_ERAM_SKIP                        ("False"),
		.IS_COMPRESSED_IMAGE                 ("False")
	) onchip_flash_0 (
		.clock                   (altpll_0_c0_clk),                                     //    clk.clk
		.reset_n                 (~rst_controller_004_reset_out_reset),                 // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_onchip_flash_0_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_onchip_flash_0_data_read),          //       .read
		.avmm_data_writedata     (mm_interconnect_0_onchip_flash_0_data_writedata),     //       .writedata
		.avmm_data_write         (mm_interconnect_0_onchip_flash_0_data_write),         //       .write
		.avmm_data_readdata      (mm_interconnect_0_onchip_flash_0_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_onchip_flash_0_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_onchip_flash_0_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_onchip_flash_0_data_burstcount),    //       .burstcount
		.avmm_csr_addr           (mm_interconnect_0_onchip_flash_0_csr_address),        //    csr.address
		.avmm_csr_read           (mm_interconnect_0_onchip_flash_0_csr_read),           //       .read
		.avmm_csr_writedata      (mm_interconnect_0_onchip_flash_0_csr_writedata),      //       .writedata
		.avmm_csr_write          (mm_interconnect_0_onchip_flash_0_csr_write),          //       .write
		.avmm_csr_readdata       (mm_interconnect_0_onchip_flash_0_csr_readdata)        //       .readdata
	);

	Embed_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c0_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_004_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	Embed_sdram sdram (
		.clk            (altpll_0_c0_clk),                          //   clk.clk
		.reset_n        (~rst_controller_004_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (dram_addr),                                //  wire.export
		.zs_ba          (dram_ba),                                  //      .export
		.zs_cas_n       (dram_cas_n),                               //      .export
		.zs_cke         (dram_cke),                                 //      .export
		.zs_cs_n        (dram_cs_n),                                //      .export
		.zs_dq          (dram_dq),                                  //      .export
		.zs_dqm         (dram_dqm),                                 //      .export
		.zs_ras_n       (dram_ras_n),                               //      .export
		.zs_we_n        (dram_we_n)                                 //      .export
	);

	Embed_slide_pio slide_pio (
		.clk        (altpll_0_c2_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_1_slide_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_slide_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_slide_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_slide_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_slide_pio_s1_readdata),   //                    .readdata
		.in_port    (sw_export),                                 // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)              //                 irq.irq
	);

	Embed_spi_0 spi_0 (
		.clk           (altpll_0_c0_clk),                                     //              clk.clk
		.reset_n       (~rst_controller_004_reset_out_reset),                 //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver0_irq),                            //              irq.irq
		.MISO          (gsensor_MISO),                                        //         external.export
		.MOSI          (gsensor_MOSI),                                        //                 .export
		.SCLK          (gsensor_SCLK),                                        //                 .export
		.SS_n          (gsensor_SS_n)                                         //                 .export
	);

	Embed_sysid sysid (
		.clock    (altpll_0_c2_clk),                                //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	Embed_timer_0 timer_0 (
		.clk        (altpll_0_c2_clk),                         //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_1_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)        //   irq.irq
	);

	Embed_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                               //                                          altpll_0_c0.clk
		.clk_0_clk_clk                                              (clk_clk),                                                       //                                            clk_0_clk.clk
		.clk_1_clk_clk                                              (clk_0_clk),                                                     //                                            clk_1_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.master_0_clk_reset_reset_bridge_in_reset_reset             (rst_controller_001_reset_out_reset),                            //             master_0_clk_reset_reset_bridge_in_reset.reset
		.modular_adc_0_reset_sink_reset_bridge_in_reset_reset       (rst_controller_001_reset_out_reset),                            //       modular_adc_0_reset_sink_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset             (rst_controller_004_reset_out_reset),                            //             nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.master_0_master_address                                    (master_0_master_address),                                       //                                      master_0_master.address
		.master_0_master_waitrequest                                (master_0_master_waitrequest),                                   //                                                     .waitrequest
		.master_0_master_byteenable                                 (master_0_master_byteenable),                                    //                                                     .byteenable
		.master_0_master_read                                       (master_0_master_read),                                          //                                                     .read
		.master_0_master_readdata                                   (master_0_master_readdata),                                      //                                                     .readdata
		.master_0_master_readdatavalid                              (master_0_master_readdatavalid),                                 //                                                     .readdatavalid
		.master_0_master_write                                      (master_0_master_write),                                         //                                                     .write
		.master_0_master_writedata                                  (master_0_master_writedata),                                     //                                                     .writedata
		.nios2_gen2_0_data_master_address                           (nios2_gen2_0_data_master_address),                              //                             nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                          //                                                     .waitrequest
		.nios2_gen2_0_data_master_byteenable                        (nios2_gen2_0_data_master_byteenable),                           //                                                     .byteenable
		.nios2_gen2_0_data_master_read                              (nios2_gen2_0_data_master_read),                                 //                                                     .read
		.nios2_gen2_0_data_master_readdata                          (nios2_gen2_0_data_master_readdata),                             //                                                     .readdata
		.nios2_gen2_0_data_master_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                        //                                                     .readdatavalid
		.nios2_gen2_0_data_master_write                             (nios2_gen2_0_data_master_write),                                //                                                     .write
		.nios2_gen2_0_data_master_writedata                         (nios2_gen2_0_data_master_writedata),                            //                                                     .writedata
		.nios2_gen2_0_data_master_debugaccess                       (nios2_gen2_0_data_master_debugaccess),                          //                                                     .debugaccess
		.nios2_gen2_0_instruction_master_address                    (nios2_gen2_0_instruction_master_address),                       //                      nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                (nios2_gen2_0_instruction_master_waitrequest),                   //                                                     .waitrequest
		.nios2_gen2_0_instruction_master_read                       (nios2_gen2_0_instruction_master_read),                          //                                                     .read
		.nios2_gen2_0_instruction_master_readdata                   (nios2_gen2_0_instruction_master_readdata),                      //                                                     .readdata
		.nios2_gen2_0_instruction_master_readdatavalid              (nios2_gen2_0_instruction_master_readdatavalid),                 //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                  //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                    //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                     //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                 //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),                //                                                     .writedata
		.altpll_1_pll_slave_address                                 (mm_interconnect_0_altpll_1_pll_slave_address),                  //                                   altpll_1_pll_slave.address
		.altpll_1_pll_slave_write                                   (mm_interconnect_0_altpll_1_pll_slave_write),                    //                                                     .write
		.altpll_1_pll_slave_read                                    (mm_interconnect_0_altpll_1_pll_slave_read),                     //                                                     .read
		.altpll_1_pll_slave_readdata                                (mm_interconnect_0_altpll_1_pll_slave_readdata),                 //                                                     .readdata
		.altpll_1_pll_slave_writedata                               (mm_interconnect_0_altpll_1_pll_slave_writedata),                //                                                     .writedata
		.mm_clock_crossing_bridge_0_s0_address                      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //                        mm_clock_crossing_bridge_0_s0.address
		.mm_clock_crossing_bridge_0_s0_write                        (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //                                                     .write
		.mm_clock_crossing_bridge_0_s0_read                         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //                                                     .read
		.mm_clock_crossing_bridge_0_s0_readdata                     (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //                                                     .readdata
		.mm_clock_crossing_bridge_0_s0_writedata                    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //                                                     .writedata
		.mm_clock_crossing_bridge_0_s0_burstcount                   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //                                                     .burstcount
		.mm_clock_crossing_bridge_0_s0_byteenable                   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //                                                     .byteenable
		.mm_clock_crossing_bridge_0_s0_readdatavalid                (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //                                                     .readdatavalid
		.mm_clock_crossing_bridge_0_s0_waitrequest                  (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //                                                     .waitrequest
		.mm_clock_crossing_bridge_0_s0_debugaccess                  (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //                                                     .debugaccess
		.modular_adc_0_sample_store_csr_address                     (mm_interconnect_0_modular_adc_0_sample_store_csr_address),      //                       modular_adc_0_sample_store_csr.address
		.modular_adc_0_sample_store_csr_write                       (mm_interconnect_0_modular_adc_0_sample_store_csr_write),        //                                                     .write
		.modular_adc_0_sample_store_csr_read                        (mm_interconnect_0_modular_adc_0_sample_store_csr_read),         //                                                     .read
		.modular_adc_0_sample_store_csr_readdata                    (mm_interconnect_0_modular_adc_0_sample_store_csr_readdata),     //                                                     .readdata
		.modular_adc_0_sample_store_csr_writedata                   (mm_interconnect_0_modular_adc_0_sample_store_csr_writedata),    //                                                     .writedata
		.modular_adc_0_sequencer_csr_address                        (mm_interconnect_0_modular_adc_0_sequencer_csr_address),         //                          modular_adc_0_sequencer_csr.address
		.modular_adc_0_sequencer_csr_write                          (mm_interconnect_0_modular_adc_0_sequencer_csr_write),           //                                                     .write
		.modular_adc_0_sequencer_csr_read                           (mm_interconnect_0_modular_adc_0_sequencer_csr_read),            //                                                     .read
		.modular_adc_0_sequencer_csr_readdata                       (mm_interconnect_0_modular_adc_0_sequencer_csr_readdata),        //                                                     .readdata
		.modular_adc_0_sequencer_csr_writedata                      (mm_interconnect_0_modular_adc_0_sequencer_csr_writedata),       //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_address                       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),        //                         nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),          //                                                     .write
		.nios2_gen2_0_debug_mem_slave_read                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),           //                                                     .read
		.nios2_gen2_0_debug_mem_slave_readdata                      (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),       //                                                     .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                     (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),      //                                                     .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                    (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),     //                                                     .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),    //                                                     .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                   (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),    //                                                     .debugaccess
		.onchip_flash_0_csr_address                                 (mm_interconnect_0_onchip_flash_0_csr_address),                  //                                   onchip_flash_0_csr.address
		.onchip_flash_0_csr_write                                   (mm_interconnect_0_onchip_flash_0_csr_write),                    //                                                     .write
		.onchip_flash_0_csr_read                                    (mm_interconnect_0_onchip_flash_0_csr_read),                     //                                                     .read
		.onchip_flash_0_csr_readdata                                (mm_interconnect_0_onchip_flash_0_csr_readdata),                 //                                                     .readdata
		.onchip_flash_0_csr_writedata                               (mm_interconnect_0_onchip_flash_0_csr_writedata),                //                                                     .writedata
		.onchip_flash_0_data_address                                (mm_interconnect_0_onchip_flash_0_data_address),                 //                                  onchip_flash_0_data.address
		.onchip_flash_0_data_write                                  (mm_interconnect_0_onchip_flash_0_data_write),                   //                                                     .write
		.onchip_flash_0_data_read                                   (mm_interconnect_0_onchip_flash_0_data_read),                    //                                                     .read
		.onchip_flash_0_data_readdata                               (mm_interconnect_0_onchip_flash_0_data_readdata),                //                                                     .readdata
		.onchip_flash_0_data_writedata                              (mm_interconnect_0_onchip_flash_0_data_writedata),               //                                                     .writedata
		.onchip_flash_0_data_burstcount                             (mm_interconnect_0_onchip_flash_0_data_burstcount),              //                                                     .burstcount
		.onchip_flash_0_data_readdatavalid                          (mm_interconnect_0_onchip_flash_0_data_readdatavalid),           //                                                     .readdatavalid
		.onchip_flash_0_data_waitrequest                            (mm_interconnect_0_onchip_flash_0_data_waitrequest),             //                                                     .waitrequest
		.onchip_memory2_0_s1_address                                (mm_interconnect_0_onchip_memory2_0_s1_address),                 //                                  onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                  (mm_interconnect_0_onchip_memory2_0_s1_write),                   //                                                     .write
		.onchip_memory2_0_s1_readdata                               (mm_interconnect_0_onchip_memory2_0_s1_readdata),                //                                                     .readdata
		.onchip_memory2_0_s1_writedata                              (mm_interconnect_0_onchip_memory2_0_s1_writedata),               //                                                     .writedata
		.onchip_memory2_0_s1_byteenable                             (mm_interconnect_0_onchip_memory2_0_s1_byteenable),              //                                                     .byteenable
		.onchip_memory2_0_s1_chipselect                             (mm_interconnect_0_onchip_memory2_0_s1_chipselect),              //                                                     .chipselect
		.onchip_memory2_0_s1_clken                                  (mm_interconnect_0_onchip_memory2_0_s1_clken),                   //                                                     .clken
		.sdram_s1_address                                           (mm_interconnect_0_sdram_s1_address),                            //                                             sdram_s1.address
		.sdram_s1_write                                             (mm_interconnect_0_sdram_s1_write),                              //                                                     .write
		.sdram_s1_read                                              (mm_interconnect_0_sdram_s1_read),                               //                                                     .read
		.sdram_s1_readdata                                          (mm_interconnect_0_sdram_s1_readdata),                           //                                                     .readdata
		.sdram_s1_writedata                                         (mm_interconnect_0_sdram_s1_writedata),                          //                                                     .writedata
		.sdram_s1_byteenable                                        (mm_interconnect_0_sdram_s1_byteenable),                         //                                                     .byteenable
		.sdram_s1_readdatavalid                                     (mm_interconnect_0_sdram_s1_readdatavalid),                      //                                                     .readdatavalid
		.sdram_s1_waitrequest                                       (mm_interconnect_0_sdram_s1_waitrequest),                        //                                                     .waitrequest
		.sdram_s1_chipselect                                        (mm_interconnect_0_sdram_s1_chipselect),                         //                                                     .chipselect
		.spi_0_spi_control_port_address                             (mm_interconnect_0_spi_0_spi_control_port_address),              //                               spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                               (mm_interconnect_0_spi_0_spi_control_port_write),                //                                                     .write
		.spi_0_spi_control_port_read                                (mm_interconnect_0_spi_0_spi_control_port_read),                 //                                                     .read
		.spi_0_spi_control_port_readdata                            (mm_interconnect_0_spi_0_spi_control_port_readdata),             //                                                     .readdata
		.spi_0_spi_control_port_writedata                           (mm_interconnect_0_spi_0_spi_control_port_writedata),            //                                                     .writedata
		.spi_0_spi_control_port_chipselect                          (mm_interconnect_0_spi_0_spi_control_port_chipselect)            //                                                     .chipselect
	);

	Embed_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c2_clk                                                 (altpll_0_c2_clk),                                             //                                               altpll_0_c2.clk
		.mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                          // mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_0_m0_address                           (mm_clock_crossing_bridge_0_m0_address),                       //                             mm_clock_crossing_bridge_0_m0.address
		.mm_clock_crossing_bridge_0_m0_waitrequest                       (mm_clock_crossing_bridge_0_m0_waitrequest),                   //                                                          .waitrequest
		.mm_clock_crossing_bridge_0_m0_burstcount                        (mm_clock_crossing_bridge_0_m0_burstcount),                    //                                                          .burstcount
		.mm_clock_crossing_bridge_0_m0_byteenable                        (mm_clock_crossing_bridge_0_m0_byteenable),                    //                                                          .byteenable
		.mm_clock_crossing_bridge_0_m0_read                              (mm_clock_crossing_bridge_0_m0_read),                          //                                                          .read
		.mm_clock_crossing_bridge_0_m0_readdata                          (mm_clock_crossing_bridge_0_m0_readdata),                      //                                                          .readdata
		.mm_clock_crossing_bridge_0_m0_readdatavalid                     (mm_clock_crossing_bridge_0_m0_readdatavalid),                 //                                                          .readdatavalid
		.mm_clock_crossing_bridge_0_m0_write                             (mm_clock_crossing_bridge_0_m0_write),                         //                                                          .write
		.mm_clock_crossing_bridge_0_m0_writedata                         (mm_clock_crossing_bridge_0_m0_writedata),                     //                                                          .writedata
		.mm_clock_crossing_bridge_0_m0_debugaccess                       (mm_clock_crossing_bridge_0_m0_debugaccess),                   //                                                          .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address                           (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                             jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                             (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),       //                                                          .write
		.jtag_uart_0_avalon_jtag_slave_read                              (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),        //                                                          .read
		.jtag_uart_0_avalon_jtag_slave_readdata                          (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                          .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                         (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                          .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                       (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                          .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                        (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                          .chipselect
		.led_pio_s1_address                                              (mm_interconnect_1_led_pio_s1_address),                        //                                                led_pio_s1.address
		.led_pio_s1_write                                                (mm_interconnect_1_led_pio_s1_write),                          //                                                          .write
		.led_pio_s1_readdata                                             (mm_interconnect_1_led_pio_s1_readdata),                       //                                                          .readdata
		.led_pio_s1_writedata                                            (mm_interconnect_1_led_pio_s1_writedata),                      //                                                          .writedata
		.led_pio_s1_chipselect                                           (mm_interconnect_1_led_pio_s1_chipselect),                     //                                                          .chipselect
		.slide_pio_s1_address                                            (mm_interconnect_1_slide_pio_s1_address),                      //                                              slide_pio_s1.address
		.slide_pio_s1_write                                              (mm_interconnect_1_slide_pio_s1_write),                        //                                                          .write
		.slide_pio_s1_readdata                                           (mm_interconnect_1_slide_pio_s1_readdata),                     //                                                          .readdata
		.slide_pio_s1_writedata                                          (mm_interconnect_1_slide_pio_s1_writedata),                    //                                                          .writedata
		.slide_pio_s1_chipselect                                         (mm_interconnect_1_slide_pio_s1_chipselect),                   //                                                          .chipselect
		.sysid_control_slave_address                                     (mm_interconnect_1_sysid_control_slave_address),               //                                       sysid_control_slave.address
		.sysid_control_slave_readdata                                    (mm_interconnect_1_sysid_control_slave_readdata),              //                                                          .readdata
		.timer_0_s1_address                                              (mm_interconnect_1_timer_0_s1_address),                        //                                                timer_0_s1.address
		.timer_0_s1_write                                                (mm_interconnect_1_timer_0_s1_write),                          //                                                          .write
		.timer_0_s1_readdata                                             (mm_interconnect_1_timer_0_s1_readdata),                       //                                                          .readdata
		.timer_0_s1_writedata                                            (mm_interconnect_1_timer_0_s1_writedata),                      //                                                          .writedata
		.timer_0_s1_chipselect                                           (mm_interconnect_1_timer_0_s1_chipselect)                      //                                                          .chipselect
	);

	Embed_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c2_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_0_c2_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (altpll_0_c2_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_0_clk),                          //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~reset_0_reset_n),                       // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_0_reset_n),                       // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (clk_0_clk),                              //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~reset_0_reset_n),                       // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (altpll_0_c2_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_0_reset_n),                       // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (),                                       //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~reset_0_reset_n),                       // reset_in1.reset
		.reset_in2      (nios2_gen2_0_debug_reset_request_reset), // reset_in2.reset
		.reset_in3      (master_0_master_reset_reset),            // reset_in3.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
